------------------------------------------------------------------
-- Company:
-- Engineer:
-- 
-- Create Date: ${DATE}
-- Design Name: 
-- Module Name: ${MODULE} - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision: 
-- Additional Comments: 
-- 
------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
--library UNISIM;
--use UNISIM.VComponents.all;

entity aaa is
--  Port ( );
end aaa;

architecture Behavioral of aaa is

begin


end Behavioral;
