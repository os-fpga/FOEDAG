`include "def.vh"
module top(input logic a, output logic b);
   bottom bot (a, b);
   
   
endmodule // top

