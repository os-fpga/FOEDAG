`timescale 1 ps/ 1 ps 
///////////////////////////////////////////////////////////////// 
// Company: 
// Engineer: 
// Create Date: ${DATE}
// Design Name: 
// Module Name: ${MODULE}
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision: 
// Additional Comments:
// 
///////////////////////////////////////////////////////////////// 


module ${MODULE}( 

    ); 
endmodule 
