module top (input logic [1:0] a, output logic [1:0] b);
assign b = a;
endmodule
